`timescale 1ns / 1ps

module instr_mem (
    input  logic [31:0] instr_rAddr,
    output logic [31:0] instr_code
);
    logic [31:0] rom [0:63];

    initial begin

        //for (int i = 0; i < 64; i++) begin
        //    rom[i] = 32'hffff_0000 + i;
        //end

        rom [0] = 32'h00000000;

        // R-Type
        //rom [1] = 32'h00208ab3; // add  x21, x1, x2
        //rom [2] = 32'h40418ab3; // sub  x21, x3, x4
        //rom [3] = 32'h00629ab3; // sll  x21, x5, x6
        //rom [4] = 32'h0083dab3; // srl  x21, x7, x8
        //rom [5] = 32'h40a4dab3; // sra  x21, x9, x10
        //rom [6] = 32'h00c5aab3; // slt  x21, x11, x12
        //rom [7] = 32'h00e6bab3; // sltu x21, x13, x14
        //rom [8] = 32'h0107cab3; // xor  x21, x15, x16
        //rom [9] = 32'h0128eab3; // or   x21, x17, x18
        //rom [10] = 32'h0149fab3; // and  x21, x19, x20

        // ADD  : 3 + 5 = 8
        // SUB  : 0 - 1 = -1
        // SLL  : 8 << 2 = 32
        // SRL  : 8 >> 2 = 2
        // SRA  : -16 >>> 4 = -1
        // SLT  : -1 < 1 = True
        // SLTU : -1(4294967295) < 1 = False
        // XOR  : 110 ^ 011 = 101(5)
        // OR   : 110 | 011 = 111(7)
        // AND  : 110 ^ 011 = 010(2)

        // S-Type
        //rom [1] = 32'h019b00a3; // sb x25, 1(x22)
        //rom [2] = 32'h019b9123; // sh x25, 2(x23)
        //rom [3] = 32'h019c2023; // sw x25, 0(x24)

        // IL-Type
        rom [1] = 32'b000000001100_00001_000_00101_0000011; // lb  x5, 12(x1)
        rom [2] = 32'b000000001100_00010_001_00101_0000011; // lh  x5, 12(x2)
        rom [3] = 32'b000000001100_00000_010_00101_0000011; // lw  x5, 12(x0)
        rom [4] = 32'b000000001100_00000_100_00101_0000011; // lbu x5, 12(x0)
        rom [5] = 32'b000000001100_00000_101_00101_0000011; // lhu x5, 12(x0)

        // IR-Type (x6 = "6" / x7 = "4294967280(-16)")
        //rom [1] = 32'b000000010000_00110_000_01000_0010011;  // addi  x8, x6, 16  (rd = rs1 + 16)
        //rom [2] = 32'b000000010000_00111_010_01000_0010011;  // slti  x8, x7, 16  (rd = rs1 < 16)
        //rom [3] = 32'b000000010000_00111_011_01000_0010011;  // sltiu x8, x7, 16  (rd = rs1 < 16)
        //rom [4] = 32'b000000010000_00110_100_01000_0010011;  // xori  x8, x6, 16  (rd = rs1 ^ 16)
        //rom [5] = 32'b000000010000_00110_110_01000_0010011;  // ori   x8, x6, 16  (rd = rs1 | 16)
        //rom [6] = 32'b000000010000_00110_111_01000_0010011;  // andi  x8, x6, 16  (rd = rs1 & 16)
        //rom [7] = 32'b0000000_00001_00110_001_01000_0010011; // slli  x8, x6, 16  (rd = rs1 << 1)
        //rom [8] = 32'b0000000_00001_00110_101_01000_0010011; // srli  x8, x6, 16  (rd = rs1 >> 1)
        //rom [9] = 32'b0100000_00100_00111_101_01000_0010011; // srai  x8, x7, 16  (rd = rs1 >>> 4)

        // B-Type
        //rom [1] = 32'b0000000_00001_00010_000_00100_1100011; // beq  x1, x2, 8 (if(rs1 == rs2) PC += imm) 
        //rom [2] = 32'b0000000_00001_00010_001_01000_1100011; // bne  x1, x2, 8 (if(rs1 != rs2) PC += imm)  
        //rom [3] = 32'b0000000_00010_00010_100_01000_1100011; // blt  x2, x2, 8 (if(rs1 <  rs2) PC += imm)  
        //rom [4] = 32'b0000000_00010_00010_101_01000_1100011; // bge  x2, x2, 8 (if(rs1 >= rs2) PC += imm)  
        //rom [5] = 32'b0000000_00010_00010_110_01000_1100011; // bltu x2, x2, 8 (if(rs1 <  rs2) PC += imm)   
        //rom [6] = 32'b0000000_00010_00010_111_01000_1100011; // bgeu x2, x2, 8 (if(rs1 >= rs2) PC += imm)

        // U-Type
        //rom [1] = 32'b00000000000000010000_00010_0110111; // lui x2, 16 (rd = imm)
        //rom [2] = 32'b00000000000000010000_00010_0010111; // aui x2, 16 (rd = PC + imm)

        // J-Type
        //rom [35] = 32'b0_0000001000_0_00000000_00010_1101111; // jal x2, 16 (rd = PC + 4, PC += imm)
        //rom [40] = 32'b000000100000_00010_000_00010_1100111;  // jalr x2, x2, 32 (rd = PC + 4, PC = rs1 + imm)
    end

    assign instr_code = rom[instr_rAddr[31:2]];

endmodule
